module somador_7b(
						input [5:0] in_c1, in_c2,
						output wire [6:0] out
						);

assign out = in_c1 + in_c2;
						
endmodule
