module somador(
					input[5:0] in_A, in_B,
					output wire[6:0] out);

assign out = in_A + in_B;
					
endmodule

					
