module proj1(
				 input [23:0] in,
				 input clr_n,
				 input ena_in,
				 output [23:0] out,
				 output ena_out
				 );



endmodule 